`timescale 1ns / 1ps

/******************************************************************************
 * Module: Transpose_Control_Top (WITH AUTO SCHEDULER)
 * * Description:
 * Top-level CONTROL module integrating Auto Scheduler, Main Scheduler, 
 * Address Generators, Compute FSM, and Mapper.
 * * UPDATES:
 * - Integrated Auto_Scheduler module.
 * - 'current_layer_id' and 'current_batch_id' are now OUTPUTS (status).
 * - Added 'weight_write_done' and 'ifmap_write_done' inputs for automation.
 ******************************************************************************/

module Transpose_Control_Top #(
    parameter DW         = 16,  // Data Width
    parameter NUM_BRAMS  = 16,  // Number of BRAMs
    parameter NUM_PE     = 16,  // Number of PEs
    parameter ADDR_WIDTH = 10   // Address Width
)(
    input  wire                   clk,
    input  wire                   rst_n,
    
    // ========================================================================
    // AUTOMATION INPUTS (From AXI Wrappers)
    // ========================================================================
    input  wire                   weight_write_done,
    input  wire                   ifmap_write_done,
    
    // ========================================================================
    // GLOBAL CONTROL INPUTS
    // ========================================================================
    input  wire                   ext_start,        // Manual Start Button
    input  wire [1:0]             ext_layer_id,     // Optional: Manual Layer ID set
    
    // ========================================================================
    // STATUS OUTPUTS (Generated by Auto Scheduler)
    // ========================================================================
    output wire [1:0]             current_layer_id, // Now an OUTPUT (Status)
    output wire [2:0]             current_batch_id, // Now an OUTPUT (Status)
    output wire                   scheduler_done,   // System Done
    output wire                   all_batches_done, // All batches for layer done
    output wire                   clear_output_bram,// Pulse to reset BRAM accumulators
    output wire                   auto_active,      // Debug: Auto Start Active
    
    // ========================================================================
    // OUTPUTS TO WEIGHT BRAM (Address & Enable)
    // ========================================================================
    output wire [NUM_BRAMS-1:0]            w_re,           
    output wire [NUM_BRAMS*ADDR_WIDTH-1:0] w_addr_rd_flat, 
    
    // ========================================================================
    // OUTPUTS TO IFMAP BRAM (Address & Enable)
    // ========================================================================
    output wire [NUM_BRAMS-1:0]            if_re,          
    output wire [NUM_BRAMS*ADDR_WIDTH-1:0] if_addr_rd_flat,
    output wire [3:0]                      ifmap_sel_out,  
    
    // ========================================================================
    // OUTPUTS TO SYSTOLIC ARRAY / DATA PATH (Control Signals)
    // ========================================================================
    output wire [NUM_PE-1:0]      en_weight_load,
    output wire [NUM_PE-1:0]      en_ifmap_load,
    output wire [NUM_PE-1:0]      en_psum,
    output wire [NUM_PE-1:0]      clear_psum,
    output wire [NUM_PE-1:0]      en_output,
    output wire [NUM_PE-1:0]      ifmap_sel_ctrl,
    
    // ========================================================================
    // OUTPUTS TO ACCUMULATION UNIT (Mapping Data)
    // ========================================================================
    output wire [NUM_BRAMS-1:0]    cmap_snapshot,
    output wire [NUM_BRAMS*14-1:0] omap_snapshot,
    output wire                    mapper_done_pulse
);

    // ========================================================================
    // INTERNAL WIRES (Interconnects)
    // ========================================================================

    // Auto Scheduler <-> Main Scheduler
    wire        final_start_signal;
    wire        batch_complete_signal;
    
    // Internal wires for layer/batch (connected to outputs)
    wire [1:0]  auto_layer_id;
    wire [2:0]  auto_batch_id;

    // Triggers from Scheduler to Sub-modules
    wire        start_Mapper;
    wire        start_weight;
    wire        start_ifmap;
    wire        start_transpose;

    // Config Signals
    wire [ADDR_WIDTH-1:0] if_addr_start;
    wire [ADDR_WIDTH-1:0] if_addr_end;
    wire [3:0]            ifmap_sel_in;
    wire [ADDR_WIDTH-1:0] addr_start;    
    wire [ADDR_WIDTH-1:0] addr_end;      
    wire [7:0]            Instruction_code;
    wire [8:0]            num_iterations;
    wire [8:0]            row_id;
    wire [5:0]            tile_id;
    wire [1:0]            layer_id_out_sched; // Unused, logic handled by AutoSched

    // Feedback Signals (Done to Scheduler)
    wire        done_mapper;
    wire        done_weight;
    wire        if_done;
    wire [4:0]  done_transpose;

    // Assignments to Outputs
    assign current_layer_id = auto_layer_id;
    assign current_batch_id = auto_batch_id;
    assign mapper_done_pulse = done_mapper;

    // ========================================================================
    // 1. INSTANTIATION: AUTO SCHEDULER (THE BRAIN)
    // ========================================================================
    Auto_Scheduler u_auto_sched (
        .clk                   (clk),
        .rst_n                 (rst_n),
        
        // Inputs from AXI
        .weight_write_done     (weight_write_done),
        .ifmap_write_done      (ifmap_write_done),
        
        // Manual Controls
        .ext_scheduler_start   (ext_start),
        .external_layer_id     (ext_layer_id),
        
        // Feedback from Main Scheduler
        .batch_complete_signal (batch_complete_signal),
        
        // Outputs to Main Scheduler
        .final_start_signal    (final_start_signal),
        .current_batch_id      (auto_batch_id),
        .current_layer_id      (auto_layer_id),
        
        // System Status Outputs
        .all_batches_complete  (all_batches_done),
        .layer_transition      (), // Internal use / debug
        .clear_output_bram     (clear_output_bram),
        .auto_start_active     (auto_active),
        .data_load_ready       ()
    );

    // ========================================================================
    // 2. INSTANTIATION: MAIN SCHEDULER_FSM
    // ========================================================================
    Scheduler_FSM #(
        .ADDR_WIDTH(ADDR_WIDTH)
    ) u_scheduler (
        .clk              (clk),
        .rst_n            (rst_n),
        .start            (final_start_signal), // Driven by Auto Scheduler
        
        // Config Inputs (Driven by Auto Scheduler)
        .current_layer_id (auto_layer_id),
        .current_batch_id (auto_batch_id),
        
        // Feedback Inputs
        .done_mapper      (done_mapper),
        .done_weight      (done_weight),
        .if_done          (if_done),
        .done_transpose   (done_transpose),
        
        // Trigger Outputs
        .start_Mapper     (start_Mapper),
        .start_weight     (start_weight),
        .start_ifmap      (start_ifmap),
        .start_transpose  (start_transpose),
        
        // Config Outputs
        .if_addr_start    (if_addr_start),
        .if_addr_end      (if_addr_end),
        .ifmap_sel_in     (ifmap_sel_in),
        .addr_start       (addr_start),
        .addr_end         (addr_end),
        .Instruction_code_transpose (Instruction_code),
        .num_iterations   (num_iterations),
        .row_id           (row_id),
        .tile_id          (tile_id),
        .layer_id         (layer_id_out_sched),
        
        // Status Outputs
        .done             (scheduler_done),
        .batch_complete   (batch_complete_signal) // Feedback loop to Auto Sched
    );

    // ========================================================================
    // 3. INSTANTIATION: COUNTER WEIGHT
    // ========================================================================
    Counter_Weight_BRAM #(
        .NUM_BRAMS  (NUM_BRAMS),
        .ADDR_WIDTH (ADDR_WIDTH)
    ) u_counter_weight (
        .clk        (clk),
        .rst_n      (rst_n),
        .start      (start_weight),     
        .addr_start (addr_start),       
        .addr_end   (addr_end),         
        
        .w_re       (w_re),             
        .w_addr_rd_flat (w_addr_rd_flat), 
        .done       (done_weight)       
    );

    // ========================================================================
    // 4. INSTANTIATION: COUNTER IFMAP
    // ========================================================================
    Counter_Ifmap_BRAM #(
        .NUM_BRAMS  (NUM_BRAMS),
        .ADDR_WIDTH (ADDR_WIDTH)
    ) u_counter_ifmap (
        .clk           (clk),
        .rst_n         (rst_n),
        .start         (start_ifmap),    
        .if_addr_start (if_addr_start),  
        .if_addr_end   (if_addr_end),    
        .ifmap_sel_in  (ifmap_sel_in),   
        
        .if_re         (if_re),            
        .if_addr_rd_flat (if_addr_rd_flat), 
        .ifmap_sel_out (ifmap_sel_out),    
        .if_done       (if_done)           
    );

    // ========================================================================
    // 5. INSTANTIATION: TRANSPOSE MATRIX FSM (COMPUTE CONTROL)
    // ========================================================================
    Transpose_Matrix_FSM #(
        .DW     (DW),
        .NUM_PE (NUM_PE)
    ) u_transpose_fsm (
        .clk              (clk),
        .rst_n            (rst_n),
        .start            (start_transpose),  
        .Instruction_code (Instruction_code), 
        .num_iterations   (num_iterations),   
        
        .en_weight_load   (en_weight_load),
        .en_ifmap_load    (en_ifmap_load),
        .en_psum          (en_psum),
        .clear_psum       (clear_psum),
        .en_output        (en_output),
        .ifmap_sel_ctrl   (ifmap_sel_ctrl),
        
        .done             (done_transpose),   
        .iter_count       ()                  
    );

    // ========================================================================
    // 6. INSTANTIATION: MM2IM MAPPER
    // ========================================================================
    MM2IM_Top #(
        .NUM_PE (NUM_PE)
    ) u_mm2im (
        .clk           (clk),
        .rst_n         (rst_n),
        .start         (start_Mapper),    
        
        .row_id        (row_id),
        .tile_id       (tile_id),
        .layer_id      (auto_layer_id), // Use Auto Layer ID
        
        .done_PE       (done_transpose),  
        
        .cmap_snapshot (cmap_snapshot),
        .omap_snapshot (omap_snapshot),
        .done          (done_mapper)      
    );

endmodule