`timescale 1ns / 1ps

/******************************************************************************
 * Module      : Transpose_Control_Top
 * Author      : Dharma Anargya Jowandy
 * Date        : January 2026
 *
 * Description :
 * Top-level control module for the Transpose Matrix Engine.
 * Integrates the Auto-Scheduler, main Scheduler FSM, and sub-controllers
 * (weight/ifmap address generators, MM2IM mapper, and Transpose FSM) to
 * manage the complete computation flow from BRAM data loading to systolic
 * array execution.
 *
 * Functionality :
 * - Coordinates weight and input feature map (Ifmap) loading
 * - Manages automatic batch sequencing via the Auto-Scheduler
 * - Controls transpose execution and address mapping logic
 * - Generates batch completion signal for synchronization with Output Manager
 *
 * Parameters :
 * - DW         : Data width (default: 16)
 * - NUM_BRAMS  : Number of BRAM banks (default: 16)
 * - NUM_PE     : Number of processing elements (default: 16)
 * - ADDR_WIDTH : Address bus width (default: 10)
 *
 ******************************************************************************/


module Transpose_Control_Top #(
    parameter DW         = 16,
    parameter NUM_BRAMS  = 16,
    parameter NUM_PE     = 16,
    parameter ADDR_WIDTH = 10
)(
    // System Signals
    input  wire                   clk,
    input  wire                   rst_n,
    
    // Automation Inputs (From AXI Wrappers)
    input  wire                   weight_write_done,
    input  wire                   ifmap_write_done,
    
    // Global Control Inputs
    input  wire                   ext_start,
    input  wire [1:0]             ext_layer_id,
    
    // Status Outputs (Generated by Auto Scheduler)
    output wire [1:0]             current_layer_id,
    output wire [2:0]             current_batch_id,
    output wire                   scheduler_done,
    output wire                   all_batches_done,
    output wire                   clear_output_bram,
    output wire                   auto_active,
    output wire                   batch_complete_signal, // Pulse for Output Manager
    
    // Outputs to Weight BRAM
    output wire [NUM_BRAMS-1:0]            w_re,
    output wire [NUM_BRAMS*ADDR_WIDTH-1:0] w_addr_rd_flat,
    
    // Outputs to Ifmap BRAM
    output wire [NUM_BRAMS-1:0]            if_re,
    output wire [NUM_BRAMS*ADDR_WIDTH-1:0] if_addr_rd_flat,
    output wire [3:0]                      ifmap_sel_out,
    
    // Outputs to Systolic Array / Data Path
    output wire [NUM_PE-1:0]      en_weight_load,
    output wire [NUM_PE-1:0]      en_ifmap_load,
    output wire [NUM_PE-1:0]      en_psum,
    output wire [NUM_PE-1:0]      clear_psum,
    output wire [NUM_PE-1:0]      en_output,
    output wire [NUM_PE-1:0]      ifmap_sel_ctrl,
    
    // Outputs to Accumulation Unit
    output wire [NUM_BRAMS-1:0]    cmap_snapshot,
    output wire [NUM_BRAMS*14-1:0] omap_snapshot,
    output wire                    mapper_done_pulse,
    output wire [4:0]              selector_mux_transpose
);

    // ========================================================================
    // Internal Signals
    // ========================================================================
    wire        final_start_signal;
    wire        internal_batch_complete;
    
    wire [1:0]  auto_layer_id;
    wire [2:0]  auto_batch_id;

    wire        start_Mapper;
    wire        start_weight;
    wire        start_ifmap;
    wire        start_transpose;

    wire [ADDR_WIDTH-1:0] if_addr_start;
    wire [ADDR_WIDTH-1:0] if_addr_end;
    wire [3:0]            ifmap_sel_in;
    wire [ADDR_WIDTH-1:0] addr_start;
    wire [ADDR_WIDTH-1:0] addr_end;
    
    wire [7:0]            Instruction_code;
    wire [8:0]            num_iterations;
    wire [8:0]            row_id;
    wire [5:0]            tile_id;
    wire [1:0]            layer_id_out_sched;
    
    wire        done_mapper;
    wire        done_weight;
    wire        if_done;
    wire [4:0]  done_transpose;

    // ========================================================================
    // Signal Assignments
    // ========================================================================
    assign current_layer_id       = auto_layer_id;
    assign current_batch_id       = auto_batch_id;
    assign mapper_done_pulse      = done_mapper;
    assign batch_complete_signal  = internal_batch_complete; // Expose status
    assign selector_mux_transpose = done_transpose;

    // ========================================================================
    // 1. Module Instantiation: Auto Scheduler
    // ========================================================================
    Auto_Scheduler u_auto_sched (
        .clk                   (clk),
        .rst_n                 (rst_n),
        .weight_write_done     (weight_write_done),
        .ifmap_write_done      (ifmap_write_done),
        .ext_scheduler_start   (ext_start),
        .external_layer_id     (ext_layer_id),
        .batch_complete_signal (internal_batch_complete),
        .final_start_signal    (final_start_signal),
        .current_batch_id      (auto_batch_id),
        .current_layer_id      (auto_layer_id),
        .all_batches_complete  (all_batches_done),
        .layer_transition      (), // Unconnected
        .clear_output_bram     (clear_output_bram),
        .auto_start_active     (auto_active),
        .data_load_ready       ()  // Unconnected
    );

    // ========================================================================
    // 2. Module Instantiation: Main Scheduler FSM
    // ========================================================================
    Scheduler_FSM #(
        .ADDR_WIDTH(ADDR_WIDTH)
    ) u_scheduler (
        .clk              (clk),
        .rst_n            (rst_n),
        .start            (final_start_signal),
        .current_layer_id (auto_layer_id),
        .current_batch_id (auto_batch_id),
        .done_mapper      (done_mapper),
        .done_weight      (done_weight),
        .if_done          (if_done),
        .done_transpose   (done_transpose),
        
        .start_Mapper     (start_Mapper),
        .start_weight     (start_weight),
        .start_ifmap      (start_ifmap),
        .start_transpose  (start_transpose),
        
        .if_addr_start    (if_addr_start),
        .if_addr_end      (if_addr_end),
        .ifmap_sel_in     (ifmap_sel_in),
        .addr_start       (addr_start),
        .addr_end         (addr_end),
        
        .Instruction_code_transpose (Instruction_code),
        .num_iterations   (num_iterations),
        .row_id           (row_id),
        .tile_id          (tile_id),
        .layer_id         (layer_id_out_sched),
        
        .done             (scheduler_done),
        .batch_complete   (internal_batch_complete) // Internal loopback
    );

    // ========================================================================
    // 3. Module Instantiation: Weight Counter
    // ========================================================================
    Counter_Weight_BRAM #(
        .NUM_BRAMS  (NUM_BRAMS),
        .ADDR_WIDTH (ADDR_WIDTH)
    ) u_counter_weight (
        .clk            (clk),
        .rst_n          (rst_n),
        .start          (start_weight),
        .addr_start     (addr_start),
        .addr_end       (addr_end),
        .w_re           (w_re),
        .w_addr_rd_flat (w_addr_rd_flat),
        .done           (done_weight)
    );

    // ========================================================================
    // 4. Module Instantiation: Ifmap Counter
    // ========================================================================
    Counter_Ifmap_BRAM #(
        .NUM_BRAMS  (NUM_BRAMS),
        .ADDR_WIDTH (ADDR_WIDTH)
    ) u_counter_ifmap (
        .clk             (clk),
        .rst_n           (rst_n),
        .start           (start_ifmap),
        .if_addr_start   (if_addr_start),
        .if_addr_end     (if_addr_end),
        .ifmap_sel_in    (ifmap_sel_in),
        .if_re           (if_re),
        .if_addr_rd_flat (if_addr_rd_flat),
        .ifmap_sel_out   (ifmap_sel_out),
        .if_done         (if_done)
    );

    // ========================================================================
    // 5. Module Instantiation: Transpose Matrix FSM
    // ========================================================================
    Transpose_Matrix_FSM #(
        .DW     (DW),
        .NUM_PE (NUM_PE)
    ) u_transpose_fsm (
        .clk              (clk),
        .rst_n            (rst_n),
        .start            (start_transpose),
        .Instruction_code (Instruction_code),
        .num_iterations   (num_iterations),
        .en_weight_load   (en_weight_load),
        .en_ifmap_load    (en_ifmap_load),
        .en_psum          (en_psum),
        .clear_psum       (clear_psum),
        .en_output        (en_output),
        .ifmap_sel_ctrl   (ifmap_sel_ctrl),
        .done             (done_transpose),
        .iter_count       () // Unconnected
    );

    // ========================================================================
    // 6. Module Instantiation: MM2IM Mapper
    // ========================================================================
    MM2IM_Top #(
        .NUM_PE (NUM_PE)
    ) u_mm2im (
        .clk           (clk),
        .rst_n         (rst_n),
        .start         (start_Mapper),
        .row_id        (row_id),
        .tile_id       (tile_id),
        .layer_id      (auto_layer_id),
        .done_PE       (done_transpose),
        .cmap_snapshot (cmap_snapshot),
        .omap_snapshot (omap_snapshot),
        .done          (done_mapper)
    );

endmodule