module systolicarray (
    
);
endmodule